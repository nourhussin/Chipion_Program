module Receiver(
    input clk, reset, rx, s_tick,
    output reg rx_done_tick,
    output[7:0] data_out
);
    parameter DATA_BITS = 8;
    parameter STOP_BITS_TICK = 16;

    localparam idle = 2'b00;
    localparam start= 2'b01;
    localparam data = 2'b10;
    localparam stop = 2'b11;

    reg [1:0] state_reg, state_next;
    reg [3:0] s_reg, s_next;
    reg [2:0] n_reg, n_next;
    reg [7:0] b_reg, b_next;
    // Register Logic
    always @(posedge clk, posedge reset)
    begin
        if(reset)
        begin
            state_reg <= idle;
            s_reg <= 0;
            n_reg <= 0;
            b_reg <= 0;
        end

        else
        begin   
            state_reg <= state_next;
            s_reg <= s_next;
            n_reg <= n_next;
            b_reg <= b_next;
        end
    end
    // Next State Logic
    always @(*)
    begin
        state_next = state_reg;
        s_next = s_reg;
        n_next = n_reg;
        b_next = b_reg;
        rx_done_tick = 1'b0;
        case(state_reg)
            idle:
                if(~rx)
                begin
                    state_next = start;
                    s_next = 0;
                end
                

            start:
                if(s_tick)
                    if(s_reg == 7)
                    begin
                        state_next = data;
                        s_next = 0;
                        n_next = 0;
                    end
                    else
                        s_next = s_reg + 1; 

            data:
                if(s_tick)
                    if(s_reg == 15)
                    begin
                        s_next = 0;
                        b_next = {rx, b_reg[7:1]};
                        if(n_reg == DATA_BITS-1)
                            state_next = stop;
                        else
                            n_next = n_reg + 1;
                    end
                    else
                        s_next = s_reg + 1;

            stop:
                if(s_tick)
                    if(s_reg== STOP_BITS_TICK-1)
                    begin
                        state_next = idle;
                        rx_done_tick = 1'b1;
                    end
                    else
                        s_next = s_reg + 1;
        endcase
    end
    // Output Logic
    assign data_out = b_reg;
endmodule